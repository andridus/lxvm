module bif
