module etf

pub enum AllocType {
	prepared_code = 3251
}
