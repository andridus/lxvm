module main

import loader

fn main() {
	loader.start()
}
