module etf