module etf
